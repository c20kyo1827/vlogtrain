module HelloWorld;
  initial begin
    $display("Hello, wor");
  end
endmodule