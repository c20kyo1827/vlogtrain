module HelloWorld;
  initial begin
    $display("Hello, wor");
  endss
endmodule