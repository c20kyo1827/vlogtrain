module HelloWorld;
  initial begin
    $display("Hello, world!");
  end
endmodule