module HelloWorld;
  initial begin
    $display("Hello, worlddd");
  end
endmodule